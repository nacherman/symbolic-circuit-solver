* Test Resistor
R1 1 0 1k
V1 1 0 DC 1
.END
