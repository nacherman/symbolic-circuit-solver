* Comprehensive Test Netlist for make_instance
.PARAM GLOBAL_RES_VAL = 1k
.PARAM OPAMP_GAIN = 100MEG
.PARAM CAP_VAL = {0.1uF * 2}
.PARAM VSIN_AMP = 2
.PARAM VSIN_PHASE_DEG = 45

* Top Level Components
VS1 N_IN 0 DC 5V AC 10 0 SIN({0} {VSIN_AMP} {1K} {0} {0} {VSIN_PHASE_DEG}) ; Offset is 0, amp & phase from param
R_INPUT N_IN N_R_IN_OUT {GLOBAL_RES_VAL}
C_MAIN N_R_IN_OUT N_MAIN_MID {CAP_VAL}
L_MAIN N_MAIN_MID 0 1mH

* Voltage Controlled Sources
E_VCVS N_E_OUT 0 N_R_IN_OUT N_MAIN_MID {OPAMP_GAIN/1000}

* Current Controlled Sources (using VS_SENSE current)
VS_SENSE N_SENSE_IN N_SENSE_OUT DC 0V
R_SENSE_PATH N_SENSE_OUT 0 1
H_CCVS N_H_OUT 0 VS_SENSE 50
F_CCCS N_F_OUT 0 VS_SENSE 100

* Subcircuit Definition
.SUBCKT MY_RC_FILTER INPUT OUTPUT LOCAL_GND PARAM R_SUBCKT=1k C_SUBCKT=1u
R_SUB INPUT N_SUB_MID {R_SUBCKT}
C_SUB N_SUB_MID OUTPUT {C_SUBCKT}
G_VCCS_SUB OUTPUT LOCAL_GND INPUT N_SUB_MID 0.1
.ENDS MY_RC_FILTER

* Subcircuit Instantiation
X_FILTER1 N_MAIN_MID N_X_OUT 0 MY_RC_FILTER R_SUBCKT=2k C_SUBCKT={CAP_VAL/2}
R_LOAD_X N_X_OUT 0 500

.AC OMEGA 1000
.END
