* Simple DC Test for Integrated Solver
VS1 N1 0 DC 10V
R1 N1 N2 2k
R2 N2 0 3k
R3 N1 0 10k

.MEASURE DC V_N1_MEAS V(N1)
.MEASURE DC V_N2_MEAS V(N2)
.MEASURE DC I_VS1_MEAS I(VS1)
.MEASURE DC I_R1_MEAS I(R1)
.MEASURE DC P_R2_MEAS POWER(R2) ; Test power measurement

.END
